_={"a":"Sidan hittas inte","b":"Sidan du söker hittades inte.","c":"Bakåt"};